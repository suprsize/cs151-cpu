module forward_logic #(
    parameter W_SIZE = 32
) (
    input [W_SIZE-1:0] inst_fd,
    input [W_SIZE-1:0] inst_xm, 
    input [W_SIZE-1:0] inst_w,
    output AFrwd1, 
    output AFrwd2, 
    output BFrwd1, 
    output BFrwd2
);
    


endmodule
